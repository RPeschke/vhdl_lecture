


library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use work.type_conversions_pgk.all;
use work.CSV_UtilityPkg.all;



use work.registerbuffer_reader_pgk.all;


entity registerbuffer_reader_et  is
    generic (
        FileName : string := "./registerbuffer_in.csv"
    );
    port (
        clk : in std_logic ;
        data : out registerbuffer_reader_rec
    );
end entity;   

architecture Behavioral of registerbuffer_reader_et is 

  constant  NUM_COL    : integer := 3;
  signal    csv_r_data : c_integer_array(NUM_COL -1 downto 0)  := (others=>0)  ;
begin

  csv_r :entity  work.csv_read_file 
    generic map (
        FileName =>  FileName, 
        NUM_COL => NUM_COL,
        useExternalClk=>true,
        HeaderLines =>  2
    ) port map (
        clk => clk,
        Rows => csv_r_data
    );

  integer_to_slv(csv_r_data(0), data.registersin.address);
  integer_to_slv(csv_r_data(1), data.registersin.value);
  integer_to_sl(csv_r_data(2), data.registersin.clk);


end Behavioral;
    